module A(output o1, input a,b);
assign o1 = ~a | ~b; 
endmodule