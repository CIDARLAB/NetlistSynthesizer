module EspToVerilog (
in1, in2, in3, in4,
out );
input in1, in2, in3, in4;
output out;
wire w0;
assign w0 =;
assign out =  w0;
endmodule
